module seedChanger(
    
)



endmodule